CircuitMaker Text
5.6
Probes: 5
R1_2
AC Analysis
0 497 200 65280
R1_2
DC Sweep
0 497 200 65280
R1_2
Transient Analysis
0 497 200 65280
R1_2
Fourier Analysis
0 497 200 65280
R2_2
Operating Point
0 569 236 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 140 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9961490 0
0
6 Title:
5 Name:
0
0
0
7
11 Multimeter~
205 682 234 0 17 21
0 6 3 3 7 0 0 0 0 0
78 79 32 68 65 84 65 32
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
1 R
5130 0 0
2
45626.1 0
0
5 SAVE-
218 497 200 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
391 0 0
2
45626.1 0
0
7 Ground~
168 244 335 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3124 0 0
2
45626.1 0
0
9 V Source~
197 244 225 0 2 5
0 5 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3421 0 0
2
45626.1 0
0
9 Resistor~
219 467 275 0 3 5
0 2 3 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8157 0 0
2
45626.1 0
0
9 Resistor~
219 543 200 0 2 5
0 4 3
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5572 0 0
2
45626.1 0
0
9 Resistor~
219 383 200 0 2 5
0 5 4
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8901 0 0
2
45626.1 0
0
8
0 3 3 0 0 8320 0 0 1 6 0 5
567 275
567 262
724 262
724 245
710 245
3 0 3 0 0 16 0 1 0 0 2 3
710 245
707 245
710 245
0 2 3 0 0 0 0 0 1 6 0 4
568 203
624 203
624 245
654 245
0 1 2 0 0 4096 0 0 3 7 0 2
244 275
244 329
1 2 4 0 0 4224 0 6 7 0 0 2
525 200
401 200
2 2 3 0 0 128 0 5 6 0 0 4
485 275
568 275
568 200
561 200
2 1 2 0 0 8320 0 4 5 0 0 3
244 246
244 275
449 275
1 1 5 0 0 8320 0 4 7 0 0 3
244 204
244 200
365 200
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
