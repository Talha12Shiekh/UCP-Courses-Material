CircuitMaker Text
5.6
Probes: 1
R2_2
Operating Point
0 752 97 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9961490 0
0
6 Title:
5 Name:
0
0
0
10
11 Multimeter~
205 809 20 0 21 21
0 3 7 8 2 0 0 0 0 0
32 54 46 54 54 55 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM3
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
5130 0 0
2
45627.1 0
0
7 Ground~
168 692 324 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
45627.1 0
0
11 Multimeter~
205 729 18 0 21 21
0 4 9 10 3 0 0 0 0 0
32 51 46 51 51 51 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM2
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3124 0 0
2
45627.1 0
0
9 V Source~
197 693 200 0 2 5
0 4 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3421 0 0
2
45627.1 0
0
7 Ground~
168 381 247 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8157 0 0
2
45627.1 0
0
11 Multimeter~
205 567 135 0 21 21
0 5 11 12 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
45627.1 0
0
9 V Source~
197 381 143 0 2 5
0 6 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8901 0 0
2
45627.1 0
0
9 Resistor~
219 808 97 0 4 5
0 3 2 0 -1
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
45627.1 0
0
9 Resistor~
219 733 97 0 2 5
0 4 3
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4747 0 0
2
45627.1 0
0
9 Resistor~
219 490 79 0 2 5
0 6 5
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
972 0 0
2
45627.1 0
0
12
4 0 2 0 0 4096 0 1 0 0 7 4
834 43
834 82
846 82
846 97
1 0 3 0 0 4096 0 1 0 0 6 4
784 43
784 89
783 89
783 97
4 0 3 0 0 4224 0 3 0 0 6 4
754 41
754 92
755 92
755 97
0 1 4 0 0 4096 0 0 3 8 0 2
704 97
704 41
0 1 2 0 0 8192 0 0 2 7 0 3
693 260
692 260
692 318
1 2 3 0 0 144 0 8 9 0 0 2
790 97
751 97
2 2 2 0 0 8192 0 4 8 0 0 5
693 221
693 260
866 260
866 97
826 97
1 1 4 0 0 8320 0 9 4 0 0 3
715 97
693 97
693 179
0 1 2 0 0 0 0 0 5 11 0 3
385 187
381 187
381 241
1 2 5 0 0 12416 0 6 10 0 0 4
542 158
542 162
508 162
508 79
2 4 2 0 0 8320 0 7 6 0 0 4
381 164
381 187
592 187
592 158
1 1 6 0 0 4224 0 10 7 0 0 3
472 79
381 79
381 122
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
