CircuitMaker Text
5.6
Probes: 5
R1_2
AC Analysis
0 497 200 65280
R1_2
DC Sweep
0 497 200 65280
R1_2
Transient Analysis
0 497 200 65280
R1_2
Fourier Analysis
0 497 200 65280
GND
Operating Point
0 481 337 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9961490 0
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 393 347 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3178 0 0
2
45626.1 0
0
10 Capacitor~
219 359 75 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3409 0 0
2
45626.1 0
0
9 Resistor~
219 364 176 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3951 0 0
2
45626.1 0
0
9 V Source~
197 363 271 0 1 5
0 0
0
0 0 17248 90
3 10V
-11 -20 10 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8885 0 0
2
45626.1 0
0
5
1 2 0 0 0 0 0 1 4 0 0 3
393 341
393 271
384 271
2 0 0 0 0 0 0 3 0 0 3 2
382 176
451 176
2 2 0 0 0 16 0 2 4 0 0 4
368 75
451 75
451 271
384 271
1 0 0 0 0 0 0 3 0 0 5 2
346 176
267 176
1 1 0 0 0 0 0 4 2 0 0 4
342 271
267 271
267 75
350 75
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
