CircuitMaker Text
5.6
Probes: 1
r1[i]
Operating Point
0 619 202 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 20 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9961490 0
0
6 Title:
5 Name:
0
0
0
6
7 Ground~
168 479 84 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
45627.2 0
0
9 V Source~
197 509 167 0 2 5
0 6 2
0
0 0 17264 270
4 9.5V
-15 -20 13 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
391 0 0
2
45627.2 0
0
9 Resistor~
219 357 219 0 4 5
0 3 2 0 -1
0
0 0 880 90
4 1.5k
1 0 29 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3124 0 0
2
45627.2 0
0
9 Resistor~
219 423 293 0 2 5
0 3 4
0
0 0 880 0
4 1.2k
-13 -14 15 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3421 0 0
2
45627.2 0
0
9 Resistor~
219 544 291 0 2 5
0 4 5
0
0 0 880 0
4 5.6k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8157 0 0
2
45627.2 0
0
9 Resistor~
219 620 219 0 2 5
0 5 6
0
0 0 880 90
4 1.2k
1 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5572 0 0
2
45627.2 0
0
6
1 2 2 0 0 4096 0 1 2 0 0 3
479 92
479 168
487 168
2 2 2 0 0 8320 0 3 2 0 0 3
357 201
357 168
487 168
1 1 3 0 0 8320 0 4 3 0 0 3
405 293
357 293
357 237
1 2 4 0 0 4224 0 5 4 0 0 4
526 291
449 291
449 293
441 293
1 2 5 0 0 8320 0 6 5 0 0 3
620 237
620 291
562 291
1 2 6 0 0 4224 0 2 6 0 0 3
529 168
620 168
620 201
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
